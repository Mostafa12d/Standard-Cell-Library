*** SPICE deck for cell 2_cell6_sim{sch} from library project
*** Created on Mon Apr 11, 2022 12:55:39
*** Last revised on Tue Apr 12, 2022 14:04:35
*** Written on Tue Apr 12, 2022 14:04:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__2_cell6 FROM CELL 2_cell6{sch}
.SUBCKT project__2_cell6 A B C gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@14 A gnd gnd nmos-BSIM130 L=0.4U W=4.8U
Mnmos@1 net@14 B gnd gnd nmos-BSIM130 L=0.4U W=4.8U
Mnmos@2 net@18 A net@14 gnd nmos-BSIM130 L=0.4U W=4.8U
Mnmos@3 net@18 C net@14 gnd nmos-BSIM130 L=0.4U W=4.8U
Mnmos@4 OUT C net@18 gnd nmos-BSIM130 L=0.4U W=4.8U
Mnmos@5 OUT B net@18 gnd nmos-BSIM130 L=0.4U W=4.8U
Mpmos@0 net@35 C OUT vdd pmos L=0.4U W=22.4U
Mpmos@1 vdd A net@35 vdd pmos L=0.4U W=22.4U
Mpmos@2 net@37 B OUT vdd pmos L=0.4U W=22.4U
Mpmos@3 vdd A net@37 vdd pmos L=0.4U W=22.4U
Mpmos@4 net@38 C OUT vdd pmos L=0.4U W=22.4U
Mpmos@5 vdd B net@38 vdd pmos L=0.4U W=22.4U
.ENDS project__2_cell6

*** SUBCIRCUIT project__NOT FROM CELL NOT{sch}
.SUBCKT project__NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=0.8U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=5.6U
.ENDS project__NOT

.global gnd vdd

*** TOP LEVEL CELL: 2_cell6_sim{sch}
X_2_cell6@0 a b c gnd out vdd project__2_cell6
XNOT@0 gnd out NOT@0_OUT vdd project__NOT

* Spice Code nodes in cell cell '2_cell6_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 PULSE 1.8 0 0.1n 0p 0p 5n 10n
Vb b 0 DC 0
Vc c 0 DC 1.8
.trans 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(a) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(a) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
