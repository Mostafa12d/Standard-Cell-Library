*** SPICE deck for cell 2_cell5_sim{sch} from library project
*** Created on Mon Apr 11, 2022 12:55:30
*** Last revised on Tue Apr 12, 2022 14:03:58
*** Written on Tue Apr 12, 2022 14:04:07 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__2_cell5 FROM CELL 2_cell5{sch}
.SUBCKT project__2_cell5 A B C D gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT A gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mnmos@1 OUT B gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mnmos@2 OUT C net@27 gnd nmos-BSIM130 L=0.4U W=1.6U
Mnmos@3 net@27 D gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mpmos@0 net@17 C OUT vdd pmos L=0.4U W=33.6U
Mpmos@1 net@17 D OUT vdd pmos L=0.4U W=33.6U
Mpmos@2 net@39 B net@17 vdd pmos L=0.4U W=33.6U
Mpmos@3 vdd A net@39 vdd pmos L=0.4U W=33.6U
.ENDS project__2_cell5

*** SUBCIRCUIT project__NOT FROM CELL NOT{sch}
.SUBCKT project__NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=0.8U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=5.6U
.ENDS project__NOT

.global gnd vdd

*** TOP LEVEL CELL: 2_cell5_sim{sch}
X_2_cell5@1 a b c d gnd out vdd project__2_cell5
XNOT@0 gnd out NOT@0_OUT vdd project__NOT

* Spice Code nodes in cell cell '2_cell5_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 DC 0
Vb b 0 DC 0
Vc c 0 DC 1.8
Vd d 0 PULSE 1.8 0 0.1n 0p 0p 5n 10n
.trans 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(d) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(d) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
