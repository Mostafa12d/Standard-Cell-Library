*** SPICE deck for cell 2_AOI22_sim{sch} from library project
*** Created on Mon Apr 11, 2022 13:08:36
*** Last revised on Tue Apr 12, 2022 12:00:37
*** Written on Tue Apr 12, 2022 12:00:41 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__2_AOI22 FROM CELL 2_AOI22{sch}
.SUBCKT project__2_AOI22 A B C D gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@4 net@66 B gnd gnd nmos-BSIM130 L=0.8U W=3.2U
Mnmos@5 OUT A net@66 gnd nmos-BSIM130 L=0.8U W=3.2U
Mnmos@6 gnd D net@67 gnd nmos-BSIM130 L=0.8U W=3.2U
Mnmos@7 net@67 C OUT gnd nmos-BSIM130 L=0.8U W=3.2U
Mpmos@4 net@49 D OUT vdd pmos L=0.4U W=22.4U
Mpmos@5 OUT C net@49 vdd pmos L=0.4U W=22.4U
Mpmos@6 vdd A net@49 vdd pmos L=0.4U W=22.4U
Mpmos@7 net@49 B vdd vdd pmos L=0.4U W=22.4U
.ENDS project__2_AOI22

*** SUBCIRCUIT project__4_NOT FROM CELL 4_NOT{sch}
.SUBCKT project__4_NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=3.2U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=22.4U
.ENDS project__4_NOT

.global gnd vdd

*** TOP LEVEL CELL: 2_AOI22_sim{sch}
X_2_AOI22@1 a b c d gnd out vdd project__2_AOI22
X_4_NOT@0 gnd out _4_NOT@0_OUT vdd project__4_NOT

* Spice Code nodes in cell cell '2_AOI22_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 DC 1.8
Vb b 0 DC 0
Vc c 0 DC 1.8
Vd d 0 PULSE 1.8 0 0.1n 500p 500p 5n 10n
.tran 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(d) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(d) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
