*** SPICE deck for cell 2_NOR_sim{sch} from library project
*** Created on Mon Apr 11, 2022 13:34:51
*** Last revised on Tue Apr 12, 2022 13:00:07
*** Written on Tue Apr 12, 2022 13:00:15 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__2_NOR FROM CELL 2_NOR{sch}
.SUBCKT project__2_NOR A B C gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT C gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mnmos@1 OUT B gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mnmos@2 OUT A gnd gnd nmos-BSIM130 L=0.4U W=1.6U
Mpmos@3 vdd A net@67 vdd pmos L=0.4U W=33.6U
Mpmos@5 net@65 C OUT vdd pmos L=0.4U W=33.6U
Mpmos@7 net@67 B net@65 vdd pmos L=0.4U W=33.6U
.ENDS project__2_NOR

*** SUBCIRCUIT project__4_NOT FROM CELL 4_NOT{sch}
.SUBCKT project__4_NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=3.2U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=22.4U
.ENDS project__4_NOT

.global gnd vdd

*** TOP LEVEL CELL: 2_NOR_sim{sch}
X_2_NOR@0 a b c gnd out vdd project__2_NOR
X_4_NOT@0 gnd out _4_NOT@0_OUT vdd project__4_NOT

* Spice Code nodes in cell cell '2_NOR_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 DC 0
Vb b 0 DC 0
Vc c 0 PULSE 1.8 0 0.1n 500p 500p 5n 10n
.trans 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(c) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(c) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
