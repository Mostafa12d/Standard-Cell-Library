*** SPICE deck for cell AOI22_sim{sch} from library project
*** Created on Wed Apr 06, 2022 13:01:23
*** Last revised on Tue Apr 12, 2022 04:08:01
*** Written on Tue Apr 12, 2022 04:08:05 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__4_NOT FROM CELL 4_NOT{sch}
.SUBCKT project__4_NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=3.2U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=22.4U
.ENDS project__4_NOT

*** SUBCIRCUIT project__AOI22 FROM CELL AOI22{sch}
.SUBCKT project__AOI22 A B C D gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@16 B gnd gnd nmos-BSIM130 L=0.8U W=1.6U
Mnmos@1 OUT A net@16 gnd nmos-BSIM130 L=0.8U W=1.6U
Mnmos@2 gnd D net@19 gnd nmos-BSIM130 L=0.8U W=1.6U
Mnmos@3 net@19 C OUT gnd nmos-BSIM130 L=0.8U W=1.6U
Mpmos@0 net@105 D OUT vdd pmos L=0.4U W=11.2U
Mpmos@1 OUT C net@105 vdd pmos L=0.4U W=11.2U
Mpmos@2 vdd A net@105 vdd pmos L=0.4U W=11.2U
Mpmos@3 net@105 B vdd vdd pmos L=0.4U W=11.2U
.ENDS project__AOI22

.global gnd vdd

*** TOP LEVEL CELL: AOI22_sim{sch}
X_4_NOT@0 gnd out _4_NOT@0_OUT vdd project__4_NOT
XAOI22@4 a b c d gnd out vdd project__AOI22

* Spice Code nodes in cell cell 'AOI22_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 DC 1.8
Vb b 0 DC 0
Vc c 0 DC 1.8
Vd d 0 PULSE 1.8 0 0.1n 400p 400p 5n 10n
.tran 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(d) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(d) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
