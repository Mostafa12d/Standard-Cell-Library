*** SPICE deck for cell cell6_sim{sch} from library project
*** Created on Mon Apr 11, 2022 22:40:21
*** Last revised on Tue Apr 12, 2022 13:47:08
*** Written on Tue Apr 12, 2022 13:48:23 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__NOT FROM CELL NOT{sch}
.SUBCKT project__NOT gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd nmos-BSIM130 L=0.4U W=0.8U
Mpmos@0 vdd IN OUT vdd pmos L=0.4U W=5.6U
.ENDS project__NOT

*** SUBCIRCUIT project__cell6 FROM CELL cell6{sch}
.SUBCKT project__cell6 A B C gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@4 A gnd gnd nmos-BSIM130 L=0.4U W=2.4U
Mnmos@1 net@4 B gnd gnd nmos-BSIM130 L=0.4U W=2.4U
Mnmos@2 net@19 A net@4 gnd nmos-BSIM130 L=0.4U W=2.4U
Mnmos@3 net@19 C net@4 gnd nmos-BSIM130 L=0.4U W=2.4U
Mnmos@4 OUT C net@19 gnd nmos-BSIM130 L=0.4U W=2.4U
Mnmos@5 OUT B net@19 gnd nmos-BSIM130 L=0.4U W=2.4U
Mpmos@0 net@39 C OUT vdd pmos L=0.4U W=11.2U
Mpmos@1 vdd A net@39 vdd pmos L=0.4U W=11.2U
Mpmos@2 net@40 B OUT vdd pmos L=0.4U W=11.2U
Mpmos@3 vdd A net@40 vdd pmos L=0.4U W=11.2U
Mpmos@4 net@41 C OUT vdd pmos L=0.4U W=11.2U
Mpmos@5 vdd B net@41 vdd pmos L=0.4U W=11.2U
.ENDS project__cell6

.global gnd vdd

*** TOP LEVEL CELL: cell6_sim{sch}
XNOT@1 gnd out NOT@1_OUT vdd project__NOT
Xcell6@0 a b c gnd out vdd project__cell6

* Spice Code nodes in cell cell 'cell6_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 PULSE 1.8 0 0.1n 0p 0p 5n 10n
Vb b 0 DC 0
Vc c 0 DC 1.8
.trans 0 100n
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(a) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(a) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
