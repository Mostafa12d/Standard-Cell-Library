*** SPICE deck for cell 2_cell7_sim{sch} from library project
*** Created on Tue Apr 12, 2022 12:08:52
*** Last revised on Tue Apr 12, 2022 12:10:10
*** Written on Tue Apr 12, 2022 12:10:22 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project__2_cell7 FROM CELL 2_cell7{sch}
.SUBCKT project__2_cell7 A B C D gnd OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 C gnd gnd nmos-BSIM130 L=0.4U W=3.2U
Mnmos@1 OUT A net@0 gnd nmos-BSIM130 L=0.4U W=3.2U
Mnmos@2 OUT A net@7 gnd nmos-BSIM130 L=0.4U W=3.2U
Mnmos@3 OUT B net@7 gnd nmos-BSIM130 L=0.4U W=3.2U
Mnmos@4 OUT C net@7 gnd nmos-BSIM130 L=0.4U W=3.2U
Mnmos@5 net@7 D gnd gnd nmos-BSIM130 L=0.4U W=3.2U
Mpmos@0 net@27 C OUT vdd pmos L=0.4U W=44.8U
Mpmos@1 net@26 B net@27 vdd pmos L=0.4U W=44.8U
Mpmos@2 net@23 A net@26 vdd pmos L=0.4U W=44.8U
Mpmos@3 net@23 D OUT vdd pmos L=0.4U W=44.8U
Mpmos@4 vdd A net@23 vdd pmos L=0.4U W=44.8U
Mpmos@5 vdd C net@23 vdd pmos L=0.4U W=44.8U
.ENDS project__2_cell7

.global gnd vdd

*** TOP LEVEL CELL: 2_cell7_sim{sch}
X_2_cell7@0 a b c d gnd out vdd project__2_cell7

* Spice Code nodes in cell cell '2_cell7_sim{sch}'
Vdd VDD 0 DC 1.8
Vgnd GND 0 DC 0
Va a 0 DC 1.8
Vb b 0 DC 0
Vc c 0 DC 0
Vd d 0 PULSE 1.8 0 0.1n 0p 0p 5n 10n
.tran 0 100n
cload out 0 9fF
.measure tran tf trig v(out) val=1.62 fall=1 TARG v(out) val=0.18 fall=1
.measure tpdr v(d) val=0.9 fall=1 TARG v(out) val=0.9 rise=1
.measure tpdf v(d) val=0.9 rise=1 TARG v(out) val=0.9 fall=1
.measure trise trig v(out) val=0.18 rise=1 TARG v(out) val=1.62 rise=1
.include "D:\University\Spring 2022\DD2\Project\BSIMTransistorModel.txt"
.END
